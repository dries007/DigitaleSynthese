-- typedef segments

package pkg_segments is
    type segment is (SEG_A, SEG_B, SEG_C, SEG_D, SEG_E);
end package;
