-- Dries Kennes
-- Datalayer
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity datalayer is
    port (
        clk: in std_logic;
        clk_en: in std_logic;
        rst: in std_logic
        -- todo  
    );
end entity;

architecture structural of datalayer is
    -- todo

begin
    -- todo

end architecture;
